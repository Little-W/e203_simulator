`ifndef DEFINE_SVH
`define DEFINE_SVH
`define SA_SIZE 16
`define ICB_LEN_W $clog2(`SA_SIZE)
`endif
